library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.conv_std_logic_vector;
use ieee.std_logic_unsigned.all;

entity tx_data is 
	PORT
	(
		signal clk16m : in std_logic;
		signal reset_n : in std_logic;
		signal next_sym_en : in std_logic;
		signal tx_data_sym : out std_logic_vector(31 downto 0)
	);
end tx_data;

architecture rtl of tx_data is

signal outdata_reg : std_logic_vector(31 downto 0);

begin

	tx_data_sym <= outdata_reg;
   set_p16m : process (clk16m)
   begin
		if (rising_edge(clk16m)) then
			if (reset_n = '0') then
				outdata_reg <= (others => '0');
			else
				if (next_sym_en = '1') then
					if (conv_integer(outdata_reg) > 128) then
						outdata_reg <= (others => '0');
					else
						outdata_reg <= outdata_reg + 1;
					end if;
				end if;
			end if;
		end if;
	end process;

--   set_p16m : process (clk16m)
--	variable cnt1 : std_logic_vector (16 downto 0);
--   begin
--		if (rising_edge(clk16m)) then
--			if (reset_n = '0') then
--				cnt1 := (others => '0');
--				outdata_reg <= (others => '0');
--			else
--				cnt1 := cnt1 + 1;
--				if (cnt1 = 0) then
--					if (conv_integer(outdata_reg) < 128) then
--						outdata_reg <= outdata_reg + 1;
--					else
--						outdata_reg <= (others => '0');
--					end if;
--				end if;
--			end if;
--		end if;
--	end process;

end rtl;
